interface intf(input logic clk,rst);
logic [1:0]ctrl;
logic [7:0]d;
logic [7:0]q;
endinterface
