`include "transaction.sv"
`include "generator.sv"
`include "intf.sv"
`include "driver.sv"
`include "environment.sv"


`include "test.sv"


`include "top.sv"
`include "usr.v"



